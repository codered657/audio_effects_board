library ieee;
use ieee.std_logic_1164.all;

use work.GeneralFuncPkg.all;

package AC97ControllerPkg is
    constant DEBUG_SINE : slv_20_vector(0 to 100) := (
        "01111101011000110100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111101011000110100",
        "01111101100010000100",
        "01111101011000110100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111111111111111100",
        "01111111110110101100",
        "01111111111111111100",
        "01111101100010000100",
        "01111101011000110100"
    );
    constant DEBUG_SQUARE : slv_20_vector(0 to 100) := (
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "01111111111111111111",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000",
        "00000000000000000000"
    );    
end package AC97ControllerPkg;



